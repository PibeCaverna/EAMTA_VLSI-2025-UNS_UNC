magic
tech sky130A
magscale 1 2
timestamp 1742412190
<< poly >>
rect 180 552 210 570
rect 268 552 298 594
rect 180 520 298 552
rect 268 268 298 520
rect 356 550 386 594
rect 444 550 474 568
rect 356 518 474 550
rect 356 262 386 518
<< metal1 >>
rect 224 860 256 1008
rect 292 982 352 1036
rect 312 918 520 948
rect 312 866 344 918
rect 488 868 520 918
rect 134 552 168 602
rect 310 552 344 604
rect 132 522 344 552
rect 398 504 432 592
rect 398 482 480 504
rect 400 474 480 482
rect 0 408 398 440
rect 448 412 480 474
rect 0 406 360 408
rect 448 370 640 412
rect 0 310 230 346
rect 448 320 480 370
rect 310 286 480 320
rect 310 234 344 286
rect 222 220 254 232
rect 222 42 256 118
rect 224 36 256 42
rect 288 0 356 54
rect 398 42 432 118
use grid__0  grid_0 inverter
timestamp 1741966214
transform 1 0 381 0 1 8
box -61 -10 259 1053
use grid__0  grid_1
timestamp 1741966214
transform 1 0 61 0 1 10
box -61 -10 259 1053
use sky130_fd_pr__nfet_01v8_3Y5EQC  sky130_fd_pr__nfet_01v8_3Y5EQC_0 inverter
timestamp 1647014411
transform 1 0 373 0 1 324
box -39 66 39 132
use sky130_fd_pr__nfet_01v8_KRUHEH__0  sky130_fd_pr__nfet_01v8_KRUHEH_0
timestamp 1741747310
transform 1 0 283 0 1 175
box -73 -101 73 101
use sky130_fd_pr__nfet_01v8_KRUHEH__0  sky130_fd_pr__nfet_01v8_KRUHEH_1
timestamp 1741747310
transform 1 0 371 0 1 175
box -73 -101 73 101
use sky130_fd_pr__pfet_01v8_MDJ67A__0  sky130_fd_pr__pfet_01v8_MDJ67A_0
timestamp 1741785174
transform 1 0 459 0 1 732
box -109 -212 109 212
use sky130_fd_pr__pfet_01v8_MDJ67A__0  sky130_fd_pr__pfet_01v8_MDJ67A_2
timestamp 1741785174
transform 1 0 195 0 1 732
box -109 -212 109 212
use sky130_fd_pr__pfet_01v8_MDJ67A__0  sky130_fd_pr__pfet_01v8_MDJ67A_3
timestamp 1741785174
transform 1 0 283 0 1 732
box -109 -212 109 212
use sky130_fd_pr__pfet_01v8_MDJ67A__0  sky130_fd_pr__pfet_01v8_MDJ67A_4
timestamp 1741785174
transform 1 0 371 0 1 732
box -109 -212 109 212
use viapoly_M1  viapoly_M1_1 inverter
timestamp 1647014411
transform 1 0 168 0 1 96
box 34 198 112 264
<< labels >>
rlabel metal1 224 860 256 1008 1 vdd
rlabel poly 268 351 298 594 1 B
rlabel metal1 222 42 256 118 1 vss
rlabel poly 356 351 386 594 1 A
rlabel metal1 448 286 480 504 1 vout
<< end >>
