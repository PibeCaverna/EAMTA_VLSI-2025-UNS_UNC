magic
tech sky130A
magscale 1 2
timestamp 1742228626
<< poly >>
rect 142 567 326 597
rect -6 56 172 86
rect -6 -268 24 56
rect -6 -334 54 -268
rect 296 -283 326 567
rect 616 567 812 597
rect 616 -93 646 567
rect 468 -123 646 -93
rect 156 -313 326 -283
rect 468 -372 498 -289
rect 372 -406 498 -372
rect 168 -634 498 -604
<< metal1 >>
rect 288 982 1700 1037
rect 0 466 114 500
rect 196 466 450 500
rect 504 466 752 500
rect 840 408 1320 442
rect 960 364 1028 374
rect 1408 372 1800 414
rect 960 286 1028 296
rect 19 -92 1701 55
rect 116 -406 338 -372
rect 1002 -391 1012 -339
rect 1064 -391 1074 -339
rect 520 -449 832 -407
rect 287 -1071 1693 -1021
<< via1 >>
rect 960 296 1028 364
rect 1012 -391 1064 -339
<< metal2 >>
rect 0 296 960 364
rect 1028 296 1038 364
rect 960 -329 1028 296
rect 960 -339 1064 -329
rect 960 -391 1012 -339
rect 960 -397 1064 -391
rect 1012 -401 1064 -397
use inverter  inverter_0 /foss/designs/mag/inverter
timestamp 1742228626
transform 1 0 320 0 1 0
box 0 0 320 1063
use inverter  inverter_1
timestamp 1742228626
transform 1 0 1600 0 1 0
box 0 0 320 1063
use inverter  inverter_2
timestamp 1742228626
transform -1 0 320 0 -1 -37
box 0 0 320 1063
use NOR  NOR_0 /foss/designs/mag/NOR
timestamp 1742228626
transform 1 0 960 0 1 2
box 0 -2 640 1063
use NOR  NOR_1
timestamp 1742228626
transform -1 0 1280 0 -1 -37
box 0 -2 640 1063
use tg  tg_0 /foss/designs/mag/Tg
timestamp 1742162383
transform 1 0 0 0 1 0
box 0 0 320 1063
use tg  tg_1
timestamp 1742162383
transform 1 0 640 0 1 0
box 0 0 320 1063
use tg  tg_2
timestamp 1742162383
transform -1 0 1600 0 -1 -37
box 0 0 320 1063
use tg  tg_3
timestamp 1742162383
transform -1 0 640 0 -1 -37
box 0 0 320 1063
use viapoly_M1  viapoly_M1_0 /foss/designs/mag/inverter
timestamp 1647014411
transform 1 0 -2 0 1 -532
box 34 198 112 264
use viapoly_M1  viapoly_M1_1
timestamp 1647014411
transform 1 0 282 0 1 -620
box 34 198 112 264
<< labels >>
rlabel metal2 0 296 960 364 1 clr
rlabel space 0 466 130 500 1 D
rlabel space 1408 372 1820 414 1 vout
rlabel poly -6 -334 24 86 1 n_clk
<< end >>
