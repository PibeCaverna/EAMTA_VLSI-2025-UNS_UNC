magic
tech sky130A
magscale 1 2
timestamp 1741792786
<< nwell >>
rect 0 486 640 1063
<< nmos >>
rect 94 106 124 406
rect 182 106 212 406
rect 414 106 444 256
<< pmos >>
rect 94 620 124 920
rect 182 620 212 920
rect 414 620 444 920
<< ndiff >>
rect 36 394 94 406
rect 36 118 48 394
rect 82 118 94 394
rect 36 106 94 118
rect 124 394 182 406
rect 124 118 136 394
rect 170 118 182 394
rect 124 106 182 118
rect 212 394 270 406
rect 212 118 224 394
rect 258 118 270 394
rect 212 106 270 118
rect 356 244 414 256
rect 356 118 368 244
rect 402 118 414 244
rect 356 106 414 118
rect 444 244 502 256
rect 444 118 456 244
rect 490 118 502 244
rect 444 106 502 118
<< pdiff >>
rect 36 908 94 920
rect 36 632 48 908
rect 82 632 94 908
rect 36 620 94 632
rect 124 908 182 920
rect 124 632 136 908
rect 170 632 182 908
rect 124 620 182 632
rect 212 908 270 920
rect 212 632 224 908
rect 258 632 270 908
rect 212 620 270 632
rect 356 908 414 920
rect 356 632 368 908
rect 402 632 414 908
rect 356 620 414 632
rect 444 908 502 920
rect 444 632 456 908
rect 490 632 502 908
rect 444 620 502 632
<< ndiffc >>
rect 48 118 82 394
rect 136 118 170 394
rect 224 118 258 394
rect 368 118 402 244
rect 456 118 490 244
<< pdiffc >>
rect 48 632 82 908
rect 136 632 170 908
rect 224 632 258 908
rect 368 632 402 908
rect 456 632 490 908
<< psubdiff >>
rect 37 10 61 44
rect 261 10 285 44
rect 357 10 381 44
rect 581 10 605 44
<< nsubdiff >>
rect 36 1026 284 1027
rect 36 992 85 1026
rect 232 992 284 1026
rect 36 991 284 992
rect 356 1026 604 1027
rect 356 992 405 1026
rect 552 992 604 1026
rect 356 991 604 992
<< psubdiffcont >>
rect 61 10 261 44
rect 381 10 581 44
<< nsubdiffcont >>
rect 85 992 232 1026
rect 405 992 552 1026
<< poly >>
rect 94 920 124 946
rect 182 920 212 946
rect 414 920 444 946
rect 94 406 124 620
rect 182 406 212 620
rect 414 510 444 620
rect 340 494 406 510
rect 340 460 356 494
rect 390 460 406 494
rect 340 444 406 460
rect 414 256 444 444
rect 94 80 124 106
rect 182 80 212 106
rect 414 80 444 106
<< polycont >>
rect 356 460 390 494
<< locali >>
rect 27 1031 293 1034
rect 27 988 33 1031
rect 288 988 293 1031
rect 27 984 293 988
rect 347 1031 613 1034
rect 347 988 353 1031
rect 608 988 613 1031
rect 347 984 613 988
rect 48 908 82 924
rect 48 616 82 632
rect 136 908 170 924
rect 136 616 170 632
rect 224 908 258 924
rect 224 616 258 632
rect 368 908 402 924
rect 368 616 402 632
rect 456 908 490 924
rect 456 616 490 632
rect 340 460 356 494
rect 390 460 406 494
rect 48 394 82 410
rect 48 102 82 118
rect 136 394 170 410
rect 136 102 170 118
rect 224 394 258 410
rect 224 102 258 118
rect 368 244 402 260
rect 368 102 402 118
rect 456 244 490 260
rect 456 102 490 118
<< viali >>
rect 33 1026 288 1031
rect 33 992 85 1026
rect 85 992 232 1026
rect 232 992 288 1026
rect 33 988 288 992
rect 353 1026 608 1031
rect 353 992 405 1026
rect 405 992 552 1026
rect 552 992 608 1026
rect 353 988 608 992
rect 48 632 82 908
rect 136 632 170 908
rect 224 632 258 908
rect 368 632 402 908
rect 456 632 490 908
rect 356 460 390 494
rect 48 118 82 394
rect 136 118 170 394
rect 224 118 258 394
rect 368 118 402 244
rect 456 118 490 244
rect 34 44 289 49
rect 34 10 61 44
rect 61 10 261 44
rect 261 10 289 44
rect 34 6 289 10
rect 354 44 609 49
rect 354 10 381 44
rect 381 10 581 44
rect 581 10 609 44
rect 354 6 609 10
<< metal1 >>
rect 21 1031 300 1037
rect 21 988 33 1031
rect 288 988 300 1031
rect 21 982 300 988
rect 341 1031 620 1037
rect 341 988 353 1031
rect 608 988 620 1031
rect 341 982 620 988
rect 42 908 88 982
rect 42 632 48 908
rect 82 632 88 908
rect 42 620 88 632
rect 130 908 176 920
rect 130 632 136 908
rect 170 632 176 908
rect 130 500 176 632
rect 218 908 264 982
rect 218 632 224 908
rect 258 632 264 908
rect 218 620 264 632
rect 362 908 408 982
rect 362 632 368 908
rect 402 632 408 908
rect 362 620 408 632
rect 450 908 496 920
rect 450 632 456 908
rect 490 632 496 908
rect 130 494 402 500
rect 130 460 356 494
rect 390 460 412 494
rect 130 454 402 460
rect 130 453 176 454
rect 42 394 88 406
rect 42 118 48 394
rect 82 118 88 394
rect 42 55 88 118
rect 130 394 176 406
rect 130 118 136 394
rect 170 118 176 394
rect 130 106 176 118
rect 218 394 264 454
rect 218 118 224 394
rect 258 118 264 394
rect 218 106 264 118
rect 362 244 408 256
rect 362 118 368 244
rect 402 118 408 244
rect 362 55 408 118
rect 450 244 496 632
rect 450 118 456 244
rect 490 118 496 244
rect 450 106 496 118
rect 22 49 301 55
rect 22 6 34 49
rect 289 6 301 49
rect 22 0 301 6
rect 342 49 621 55
rect 342 6 354 49
rect 609 6 621 49
rect 342 0 621 6
<< end >>
