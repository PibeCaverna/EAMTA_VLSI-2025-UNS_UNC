magic
tech sky130A
magscale 1 2
timestamp 1741981168
<< nwell >>
rect 320 -1107 640 -530
rect 1264 -1107 1584 -530
<< nmos >>
rect 470 -294 500 -144
rect 1414 -294 1444 -144
<< pmos >>
rect 470 -978 500 -678
rect 1414 -978 1444 -678
<< ndiff >>
rect 412 -156 470 -144
rect 412 -282 424 -156
rect 458 -282 470 -156
rect 412 -294 470 -282
rect 500 -156 558 -144
rect 500 -282 512 -156
rect 546 -282 558 -156
rect 500 -294 558 -282
rect 1356 -156 1414 -144
rect 1356 -282 1368 -156
rect 1402 -282 1414 -156
rect 1356 -294 1414 -282
rect 1444 -156 1502 -144
rect 1444 -282 1456 -156
rect 1490 -282 1502 -156
rect 1444 -294 1502 -282
<< pdiff >>
rect 412 -690 470 -678
rect 412 -966 424 -690
rect 458 -966 470 -690
rect 412 -978 470 -966
rect 500 -690 558 -678
rect 500 -966 512 -690
rect 546 -966 558 -690
rect 500 -978 558 -966
rect 1356 -690 1414 -678
rect 1356 -966 1368 -690
rect 1402 -966 1414 -690
rect 1356 -978 1414 -966
rect 1444 -690 1502 -678
rect 1444 -966 1456 -690
rect 1490 -966 1502 -690
rect 1444 -978 1502 -966
<< ndiffc >>
rect 424 -282 458 -156
rect 512 -282 546 -156
rect 1368 -282 1402 -156
rect 1456 -282 1490 -156
<< pdiffc >>
rect 424 -966 458 -690
rect 512 -966 546 -690
rect 1368 -966 1402 -690
rect 1456 -966 1490 -690
<< psubdiff >>
rect 355 -88 379 -54
rect 579 -88 603 -54
rect 1299 -88 1323 -54
rect 1523 -88 1547 -54
<< nsubdiff >>
rect 356 -1036 604 -1035
rect 356 -1070 408 -1036
rect 555 -1070 604 -1036
rect 356 -1071 604 -1070
rect 1300 -1036 1548 -1035
rect 1300 -1070 1352 -1036
rect 1499 -1070 1548 -1036
rect 1300 -1071 1548 -1070
<< psubdiffcont >>
rect 379 -88 579 -54
rect 1323 -88 1523 -54
<< nsubdiffcont >>
rect 408 -1070 555 -1036
rect 1352 -1070 1499 -1036
<< poly >>
rect 470 -144 500 -118
rect 1414 -144 1444 -118
rect 470 -367 500 -294
rect 1414 -367 1444 -294
rect 470 -678 500 -609
rect 1414 -678 1444 -609
rect 470 -1004 500 -978
rect 1414 -1004 1444 -978
<< locali >>
rect 424 -156 458 -140
rect 424 -298 458 -282
rect 512 -156 546 -140
rect 512 -298 546 -282
rect 1368 -156 1402 -140
rect 1368 -298 1402 -282
rect 1456 -156 1490 -140
rect 1456 -298 1490 -282
rect 424 -690 458 -674
rect 424 -982 458 -966
rect 512 -690 546 -674
rect 512 -982 546 -966
rect 1368 -690 1402 -674
rect 1368 -982 1402 -966
rect 1456 -690 1490 -674
rect 1456 -982 1490 -966
rect 347 -1032 613 -1028
rect 347 -1075 352 -1032
rect 607 -1075 613 -1032
rect 347 -1078 613 -1075
rect 1291 -1032 1557 -1028
rect 1291 -1075 1296 -1032
rect 1551 -1075 1557 -1032
rect 1291 -1078 1557 -1075
<< viali >>
rect 351 -54 606 -50
rect 351 -88 379 -54
rect 379 -88 579 -54
rect 579 -88 606 -54
rect 351 -93 606 -88
rect 1295 -54 1550 -50
rect 1295 -88 1323 -54
rect 1323 -88 1523 -54
rect 1523 -88 1550 -54
rect 1295 -93 1550 -88
rect 424 -282 458 -156
rect 512 -282 546 -156
rect 1368 -282 1402 -156
rect 1456 -282 1490 -156
rect 424 -966 458 -690
rect 512 -966 546 -690
rect 1368 -966 1402 -690
rect 1456 -966 1490 -690
rect 352 -1036 607 -1032
rect 352 -1070 408 -1036
rect 408 -1070 555 -1036
rect 555 -1070 607 -1036
rect 352 -1075 607 -1070
rect 1296 -1036 1551 -1032
rect 1296 -1070 1352 -1036
rect 1352 -1070 1499 -1036
rect 1499 -1070 1551 -1036
rect 1296 -1075 1551 -1070
<< metal1 >>
rect 142 990 1728 1034
rect 142 -72 174 30
rect 178 8 460 48
rect 492 8 764 48
rect 796 8 1076 48
rect 1108 8 1394 48
rect 1426 8 1770 48
rect 339 -50 460 -44
rect 492 -50 618 -44
rect 339 -54 351 -50
rect 178 -93 351 -54
rect 606 -54 618 -50
rect 1283 -50 1394 -44
rect 1426 -50 1562 -44
rect 1283 -54 1295 -50
rect 606 -93 1295 -54
rect 1550 -93 1562 -50
rect 178 -94 1562 -93
rect 339 -99 618 -94
rect 1283 -99 1562 -94
rect 418 -156 464 -144
rect 418 -282 424 -156
rect 458 -282 464 -156
rect 418 -294 464 -282
rect 506 -156 552 -144
rect 506 -282 512 -156
rect 546 -282 552 -156
rect 506 -294 552 -282
rect 1362 -156 1408 -144
rect 1362 -282 1368 -156
rect 1402 -282 1408 -156
rect 1362 -294 1408 -282
rect 1450 -156 1496 -144
rect 1450 -282 1456 -156
rect 1490 -282 1496 -156
rect 1450 -294 1496 -282
rect 424 -678 458 -294
rect 512 -678 546 -294
rect 1368 -678 1402 -294
rect 1456 -678 1490 -294
rect 418 -690 464 -678
rect 418 -966 424 -690
rect 458 -966 464 -690
rect 418 -978 464 -966
rect 506 -690 552 -678
rect 506 -966 512 -690
rect 546 -966 552 -690
rect 506 -978 552 -966
rect 1362 -690 1408 -678
rect 1362 -966 1368 -690
rect 1402 -966 1408 -690
rect 1362 -978 1408 -966
rect 1450 -690 1496 -678
rect 1450 -966 1456 -690
rect 1490 -966 1496 -690
rect 1450 -978 1496 -966
rect 340 -1032 619 -1026
rect 340 -1034 352 -1032
rect 190 -1075 352 -1034
rect 607 -1034 619 -1032
rect 1284 -1032 1563 -1026
rect 1284 -1034 1296 -1032
rect 607 -1075 1296 -1034
rect 1551 -1075 1563 -1032
rect 190 -1076 1563 -1075
rect 340 -1081 619 -1076
rect 1284 -1081 1563 -1076
use inverter  inverter_0 /foss/designs/mag/inverter
timestamp 1741977694
transform -1 0 326 0 -1 -45
box 0 0 320 1063
use inverter  inverter_1
timestamp 1741977694
transform 1 0 1572 0 1 4
box 0 0 320 1063
use inverter  inverter_3
timestamp 1741977694
transform 1 0 312 0 1 2
box 0 0 320 1063
use NOR  NOR_0 /foss/designs/mag/NOR
timestamp 1741809433
transform 1 0 942 0 1 8
box 0 -2 640 1063
use NOR  NOR_1
timestamp 1741809433
transform -1 0 1274 0 -1 -43
box 0 -2 640 1063
use tg  tg_0 /foss/designs/mag/Tg
timestamp 1741977694
transform 1 0 626 0 1 0
box 2 2 322 1065
use tg  tg_1
timestamp 1741977694
transform 1 0 -4 0 1 2
box 2 2 322 1065
use tg  tg_2
timestamp 1741977694
transform -1 0 642 0 -1 -42
box 2 2 322 1065
use tg  tg_3
timestamp 1741977694
transform 1 0 2060 0 1 1846
box 2 2 322 1065
use tg  tg_4
timestamp 1741977694
transform -1 0 1586 0 -1 -42
box 2 2 322 1065
<< labels >>
rlabel nwell 408 -1070 555 -1036 5 vdd
rlabel poly 470 -367 500 -294 5 n_clk
rlabel poly 470 -678 500 -609 5 clk
rlabel metal1 512 -710 546 -266 5 in
rlabel metal1 424 -744 458 -268 5 out
rlabel metal1 1323 -88 1523 -54 5 vss
rlabel nwell 1352 -1070 1499 -1036 5 vdd
rlabel poly 1414 -367 1444 -294 5 n_clk
rlabel poly 1414 -678 1444 -609 5 clk
rlabel metal1 1456 -710 1490 -266 5 in
rlabel metal1 1368 -744 1402 -268 5 out
rlabel metal1 379 -88 579 -54 5 vss
<< end >>
