magic
tech sky130A
magscale 1 2
timestamp 1741785174
<< error_p >>
rect -134 156 -76 162
rect -134 122 -122 156
rect 202 137 262 175
rect 286 156 344 162
rect 286 122 298 156
rect -134 116 -76 122
rect 286 116 344 122
rect -344 -122 -286 -116
rect 76 -122 134 -116
rect -344 -156 -332 -122
rect -344 -162 -286 -156
rect -8 -175 52 -137
rect 76 -156 88 -122
rect 76 -162 134 -156
<< nwell >>
rect -218 137 8 175
rect 202 137 428 175
rect -428 -137 428 137
rect -428 -175 -202 -137
rect -8 -175 218 -137
<< pmos >>
rect -330 -75 -300 75
rect -120 -75 -90 75
rect 90 -75 120 75
rect 300 -75 330 75
<< pdiff >>
rect -392 63 -330 75
rect -392 -63 -380 63
rect -346 -63 -330 63
rect -392 -75 -330 -63
rect -300 63 -238 75
rect -300 -63 -284 63
rect -250 -63 -238 63
rect -300 -75 -238 -63
rect -182 63 -120 75
rect -182 -63 -170 63
rect -136 -63 -120 63
rect -182 -75 -120 -63
rect -90 63 -28 75
rect -90 -63 -74 63
rect -40 -63 -28 63
rect -90 -75 -28 -63
rect 28 63 90 75
rect 28 -63 40 63
rect 74 -63 90 63
rect 28 -75 90 -63
rect 120 63 182 75
rect 120 -63 136 63
rect 170 -63 182 63
rect 120 -75 182 -63
rect 238 63 300 75
rect 238 -63 250 63
rect 284 -63 300 63
rect 238 -75 300 -63
rect 330 63 392 75
rect 330 -63 346 63
rect 380 -63 392 63
rect 330 -75 392 -63
<< pdiffc >>
rect -380 -63 -346 63
rect -284 -63 -250 63
rect -170 -63 -136 63
rect -74 -63 -40 63
rect 40 -63 74 63
rect 136 -63 170 63
rect 250 -63 284 63
rect 346 -63 380 63
<< poly >>
rect -138 156 -72 172
rect -138 122 -122 156
rect -88 122 -72 156
rect -138 106 -72 122
rect 282 156 348 172
rect 282 122 298 156
rect 332 122 348 156
rect 282 106 348 122
rect -330 75 -300 101
rect -120 75 -90 106
rect 90 75 120 101
rect 300 75 330 106
rect -330 -106 -300 -75
rect -120 -101 -90 -75
rect 90 -106 120 -75
rect 300 -101 330 -75
rect -348 -122 -282 -106
rect -348 -156 -332 -122
rect -298 -156 -282 -122
rect -348 -172 -282 -156
rect 72 -122 138 -106
rect 72 -156 88 -122
rect 122 -156 138 -122
rect 72 -172 138 -156
<< polycont >>
rect -122 122 -88 156
rect 298 122 332 156
rect -332 -156 -298 -122
rect 88 -156 122 -122
<< locali >>
rect -138 122 -122 156
rect -88 122 -72 156
rect 282 122 298 156
rect 332 122 348 156
rect -380 63 -346 79
rect -380 -79 -346 -63
rect -284 63 -250 79
rect -284 -79 -250 -63
rect -170 63 -136 79
rect -170 -79 -136 -63
rect -74 63 -40 79
rect -74 -79 -40 -63
rect 40 63 74 79
rect 40 -79 74 -63
rect 136 63 170 79
rect 136 -79 170 -63
rect 250 63 284 79
rect 250 -79 284 -63
rect 346 63 380 79
rect 346 -79 380 -63
rect -348 -156 -332 -122
rect -298 -156 -282 -122
rect 72 -156 88 -122
rect 122 -156 138 -122
<< viali >>
rect -122 122 -88 156
rect 298 122 332 156
rect -380 -63 -346 63
rect -284 -63 -250 63
rect -170 -63 -136 63
rect -74 -63 -40 63
rect 40 -63 74 63
rect 136 -63 170 63
rect 250 -63 284 63
rect 346 -63 380 63
rect -332 -156 -298 -122
rect 88 -156 122 -122
<< metal1 >>
rect -134 156 -76 162
rect -134 122 -122 156
rect -88 122 -76 156
rect -134 116 -76 122
rect 286 156 344 162
rect 286 122 298 156
rect 332 122 344 156
rect 286 116 344 122
rect -386 63 -340 75
rect -386 -63 -380 63
rect -346 -63 -340 63
rect -386 -75 -340 -63
rect -290 63 -244 75
rect -290 -63 -284 63
rect -250 -63 -244 63
rect -290 -75 -244 -63
rect -176 63 -130 75
rect -176 -63 -170 63
rect -136 -63 -130 63
rect -176 -75 -130 -63
rect -80 63 -34 75
rect -80 -63 -74 63
rect -40 -63 -34 63
rect -80 -75 -34 -63
rect 34 63 80 75
rect 34 -63 40 63
rect 74 -63 80 63
rect 34 -75 80 -63
rect 130 63 176 75
rect 130 -63 136 63
rect 170 -63 176 63
rect 130 -75 176 -63
rect 244 63 290 75
rect 244 -63 250 63
rect 284 -63 290 63
rect 244 -75 290 -63
rect 340 63 386 75
rect 340 -63 346 63
rect 380 -63 386 63
rect 340 -75 386 -63
rect -344 -122 -286 -116
rect -344 -156 -332 -122
rect -298 -156 -286 -122
rect -344 -162 -286 -156
rect 76 -122 134 -116
rect 76 -156 88 -122
rect 122 -156 134 -122
rect 76 -162 134 -156
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.75 l 0.15 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
