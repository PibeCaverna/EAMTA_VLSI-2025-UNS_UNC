magic
tech sky130A
magscale 1 2
timestamp 1647014411
<< poly >>
rect -33 116 33 132
rect -33 82 -17 116
rect 17 82 33 116
rect -33 66 33 82
<< polycont >>
rect -17 82 17 116
<< locali >>
rect -33 82 -17 116
rect 17 82 33 116
<< viali >>
rect -17 82 17 116
<< metal1 >>
rect -29 116 29 122
rect -39 82 -17 116
rect 17 82 39 116
rect -29 76 29 82
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.75 l 0.150 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
